// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
// Created on Sun May 18 22:27:31 2025

// synthesis message_off 10175

`timescale 1ns/1ns

module FSM_based_traffic_controller (
    reset,clock,c,
    NS_G,NS_R,EW_G,EW_R);

    input reset;
    input clock;
    input c;
    tri0 reset;
    tri0 c;
    output NS_G;
    output NS_R;
    output EW_G;
    output EW_R;
    reg NS_G;
    reg NS_R;
    reg EW_G;
    reg EW_R;
    reg [1:0] fstate;
    reg [1:0] reg_fstate;
    parameter NS=0,EW=1;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or c)
    begin
        if (reset) begin
            reg_fstate <= NS;
            NS_G <= 1'b0;
            NS_R <= 1'b0;
            EW_G <= 1'b0;
            EW_R <= 1'b0;
        end
        else begin
            NS_G <= 1'b0;
            NS_R <= 1'b0;
            EW_G <= 1'b0;
            EW_R <= 1'b0;
            case (fstate)
                NS: begin
                    if (c)
                        reg_fstate <= EW;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= NS;

                    EW_G <= 1'b1;

                    NS_G <= 1'b0;

                    EW_R <= 1'b0;

                    NS_R <= 1'b1;
                end
                EW: begin
                    if (~(c))
                        reg_fstate <= NS;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= EW;

                    EW_G <= 1'b0;

                    NS_G <= 1'b1;

                    EW_R <= 1'b1;

                    NS_R <= 1'b0;
                end
                default: begin
                    NS_G <= 1'bx;
                    NS_R <= 1'bx;
                    EW_G <= 1'bx;
                    EW_R <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // FSM_based_traffic_controller
