module mod_7_counter_tb;

    reg clk, rst;
    wire [2:0] count;

    // Instantiate the Mod-7 counter
    mod_7_counter uut (
        .clk(clk),
        .rst(rst),
        .count(count)
    );

    // Clock Generation (50MHz, 20ns period)
    always #10 clk = ~clk;

    // Test Procedure
    initial begin
	 
        clk = 0;  
        rst = 1;  
        #20;  // Apply Reset

        rst = 0;  
        #200;  // Run for multiple clock cycles

        $finish;
    end

    // Monitor count value changes
    always @(posedge clk) begin
        $display("Time: %0t | Count: %0d", $time, count);
    end

endmodule
